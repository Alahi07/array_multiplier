// Code your design here
`include "top.v"
